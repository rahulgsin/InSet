* Version 2.0 Copyright © Linear Technology Corp. 10/19/05. All rights reserved.
*
.SUBCKT LT1192 3 nois 7 4 6 ;(+IN -IN V+ V- OUT)
* INPUT
*nois
VNoiw nois 2 dc 0 TRNOISE (2m 1n 0 0 )

RC1 7 80 11.789
RC2 7 90 11.789
Q1 80 2 10 QM1
Q2 90 3 11 QM2
CIN 2 3 1.8e-12
C1 80 90 5.5981E-11
RE1 10 12 8.6552
RE2 11 12 8.6552
IEE 12 4 0.016501
RE 12 0 12120
* INTERMEDIATE
GCM 0 8 12 0 4.7699e-6
GA 8 0 80 90 0.084823
R2 8 0 100000
C2 1 8 3e-11
GB 1 0 8 0 3.1289
RO2 1 0 1.5
* OUTPUT
RSO 1 6 1
ECL 18 0 1 6 12.252
GCL 0 8 20 0 1
RCL 20 0 10
D1 18 19 DM1
VOD1 19 20 0
D2 20 21 DM1
VOD2 21 18 0.18378
*
D3A 131 70 DM3
D3B 13 131 DM3
GPL 0 8 70 7 1
VC 13 6 2.6003
RPLA 7 70 10
RPLB 7 131 1000
D4A 60 141 DM3
D4B 141 14 DM3
GNL 0 8 60 4 1
VE 6 14 2.1003
RNLA 60 4 10
RNLB 141 4 1000
*
IP 7 4 0.015499
DSUB 4 7 DM2
* MODELS
.MODEL QM1 NPN(IS=8e-16 BF=13750)
.MODEL QM2 NPN(IS=8.0621E-16 BF=20625)
.MODEL DM1 D(IS=1e-20)
.MODEL DM2 D(IS=8e-16 BV=21.6)
.MODEL DM3 D(IS=1e-16)
.ENDS LT1192

