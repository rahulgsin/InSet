*PEAK DETECTOR SUBCIRCUIT

.include ths3001.cir
.SUBCKT PEAKDETECTOR 1 15

.MODEL germ d
+IS=1.88569e-06 RS=0.160685 N=1.03056 EG=0.634401
+XTI=0.5 BV=20 IBV=1.5e-05 CJO=1.20949e-10
+VJ=0.4 M=0.520353 FC=0.5 TT=0
+KF=0 AF=1


C1 1 2 50PF
C2 2 0 10PF
*rtemp 2 51 10k
*
*XOP1	2 3 4 5 6	LT1192
*RO1	3	0	100
*RO2	3	6	100
*CO1	6	7	15nF
*ri1	2	0	1meg
*CO2	3	0	10pf
*rl	7	0	1meg
*VCC1 	4 0 DC 15V
*VEE1	5 0 DC -15V
*

R1 2 0 100k
D1 2 8 new
C3 8 0 10pF 
R2 8 0 100k

*C3 8 0 10pF 
*R2 8 0 100k
C4 8 9 1pf
*

XOP2	9 10 11 12 13	THS3001
RO3	10	0	10
RO4	10	13	100
C03	13 	14 	1pf
ri2	9	0	1meg
*CO4	10	0	10pf
R3	14	0	10k
*rl2	13	0	75
VCC2	11 0 DC 15v
VEE2	12 0 DC -15v
*

rfilt	14	15	160
*cfilt	15	0	1pf 

.ENDS

.include lt1192.cir
XPEAK1 1 2 PEAKDETECTOR
XPEAK2 3 4 PEAKDETECTOR 

XOPdiff	5 6 7 8 9	THS3001
VCCd	7 0 DC 15v
VEEd	8 0 DC -15v

r1	2	5	10MEG
r2	4	6	10MEG
r3	5	9	10MEG
r4	6	0	10MEG

rf1	9 	10	3.3k 
rf2	10	11	3.3k
cf1	10 	0	50pf
cf2	11 	0	50pf


AVSRC1 %V([1]) filesrc1
*.include Input_signal.txt
.model filesrc1 filesource (file="dataa/x2_profilecoast_volt1.txt" )

AVSRC2 %V([3]) filesrc2
*.include Input_signal.txt
.model filesrc2 filesource (file="dataa/x1_profilecoast_volt1.txt" )

.CONTROL
*AC 	DEC 	 1k 500MEG
*PLOT mag(V(2,7)) xlog
TRAN 1ns 10us
plot v(1) v(2) v(4)
plot v(1) 
plot v(9) 
plot v(11)
*plot v(1) v(2)
*.include plotng.txt
wrdata bbqx1ext v(1)
wrdata bbqx2extd v(9) 
wrdata bbqx2ext v(11)
wrdata pick2ext v(2)
wrdata pickx2ext v(4)
*wrdata plot4 v(9)
