Cap_check

Cin 2 3 5pf
ro 3 0 100k

VIN 2 1 AC SIN(0 50m 10meg)
VCLOCK 1 0 PWL( 0 0 1US 0.2 2US 0.4 3US 0.6 4US 0.8 5US 1 6US 1.2 7US 1.4 8US 1.6 9US 1.8 10US 2 ) 
*AVSRC %V([1]) filesrc
*.model filesrc filesource (file="cap_out.data" )

.control
tran 1ns 10us
plot V(3) v(2)

