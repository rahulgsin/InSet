BUFFER

.SUBCKT buf 1 5
.include lt1192.cir
XOP	1 5 3 4 5	LT1192
VCC 	3 0 DC 15V
VEE	4 0 DC -15V
.ENDS

*Xamp 1 2 buf
*Xatt 2 3 att20
*vin 1 0 sin(0 10m 10meg)
*.control
*tran 1ns 1us
*plot v(1) V(2)
