Amplifier of 10db

.SUBCKT amp10 1 6
.include lt1192.cir
XOP	1 2 3 4 5	LT1192
R1	2	0	150
R2	2	5	500
cL	5	6	15nf
rl	6	0	10k
VCC 	3 0 DC 15V
VEE	4 0 DC -15V
.ENDS

