TOPOS SIGNAL CHAIN from BPM plates to ADC

.include att10.cir
.include att20.cir
.include att30.cir
.include amp10.cir
.include amp20.cir

*First topos chain
Rb 22 0 100k
Cb1 1 22 50pF
Cb2 22 0 50pF
*Vin 1 0 ac sin(0 1m 10meg)
AVSRC %V([1]) filesrc
*.include Input_signal.txt
.model filesrc filesource (file="daata/x1_coast_v.txt" )

*head ampliflier of 20db
*rser1	3 0 10meg
Xamp20 22 4 amp20

*second topos chain

Rb1 221 0 100k
Cb11 11 221 50pF
Cb21 221 0 50pF
*Vin1 11 0 ac sin(0 1m 10meg)
AVSRC1 %V([11]) filesrc1
*.include Input_signal.txt
.model filesrc1 filesource (file="daata/x2_coast_v.txt" )

*head ampliflier of 20db
*rser1	3 0 10meg
Xamp201 221 41 amp20

*3 tops chain

Rb11 2211 0 100k
Cb111 111 2211 50pF
Cb211 2211 0 50pF
*Vin1 111 0 ac sin(0 1m 10meg)
AVSRC11 %V([111]) filesrc11
.model filesrc11 filesource (file="daata/y1_coast_v.txt" )

Xamp2011 2211 411 amp20


*4 tops chain

Rb111 22111 0 100k
Cb1111 1111 22111 50pF
Cb2111 22111 0 50pF
*Vin1 1111 0 ac sin(0 1m 10meg)
AVSRC111 %V([1111]) filesrc111
.model filesrc111 filesource (file="daata/y2_coast_v.txt" )

Xamp20111 22111 4111 amp20


.CONTROL
*ac 	DEC 1000 1k 1000MEG
*plot db(v(4)/v(1)) xlog
*plot 180/pi*phase(V(4)/v(1)) 
tran 1ns 50us 
*plot v(1) v(11) 
*plot v(111) v(1111)
*plot v(4) v(41)
*plot v(411) v(4111)
*plot v(1) v(22) v(33) v(3)
*plot v(4)
*plot v(5)
*plot v(6)
*plot v(111) v(9)
*plot v(7) v(8) v(9) 
*.include plotng.txt
*setplot tran1
*linearize
wrdata ip v(1) 
wrdata op v(4)
*wrdata x2_coast_1 v(41)
*wrdata y1_coast_1 v(411)
*wrdata y2_coast_1 v(4111)
