
Vin 1 0 ac sin(0 100m 10meg)

OLOSSY 1 0 2 0 rg58
.model rg58 LTRA(LEN=200 R=0.048 L=0.253u G=0 C=0.101n)

Rl 2 0 50
*Y1 1 0 2 0 lossy LEN=200
*.MODEL lossy txl R=0.048 L=0.253e-6 G=0.001e-12 C=0.101e-9 length=1

*Y1 1 0 2 0 ymod LEN=2
*.MODEL ymod txl R= 0.048 L=8.972e−9 G=0 C=0.468e−12 length=16

.CONTROL
ac 	LIN 	1000 100k 100MEG
plot (vdb(2)-Vdb(1))
plot 180/pi*phase(V(2)/v(1)) 
TRAN 1NS 2US
PLOT V(1) V(2)

