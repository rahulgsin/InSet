Attenuator of -30db

.SUBCKT att30 41 11
.include lt1192.cir
XOP	0 2 3 4 5	LT1192
R1	41	2	100000
R2	2	5	3000
cL	5	6	15nf
rl	6	0	1meG
VCC 	3 0 DC 15V
VEE	4 0 DC -15V

XOPB	0 7 8 9 10	LT1192
RB1	6	7	100000
RB2	7	10	100000
cLB	10	11	15nf
rlB	11	0	1meg
VCCB 	8 0 DC 15V
VEEB	9 0 DC -15V
.ENDS

