BPM simulation program for NGspice

R1 2 0 100k

C1 1 2 50PF

C2 2 0 50PF

*vin 1 0 ac sin(0 1m 10meg)
AVSRC %V([1]) filesrc1
.model filesrc1 filesource (file="dat/x1_profile_bunched.txt" amploffset=[0 0] amplscale=[1 1]
+ timeoffset=0 timescale=1
+ timerelative=false amplstep=false)

R11 22 0 100k

C11 11 22 50PF

C21 22 0 50PF

*vin2 11 0 ac sin(0 1m 10meg)
AVSRC1 %V([11]) filesrc2
.model filesrc2 filesource (file="dat/x2_profile_bunched.txt" amploffset=[0 0] amplscale=[1 1]
+ timeoffset=0 timescale=1
+ timerelative=false amplstep=false) )

R13 23 0 100k

C13 13 23 50PF

C23 23 0 50PF

*vin3 13 0 ac sin(0 1m 10meg)
AVSRC3 %V([13]) filesrc3
.model filesrc3 filesource (file="dat/y1_profile_bunched.txt" amploffset=[0 0] amplscale=[1 1]
+ timeoffset=0 timescale=1
+ timerelative=false amplstep=false) )

R14 24 0 100k

C14 14 24 50PF

C24 24 0 50PF

*vin3 13 0 ac sin(0 1m 10meg)
AVSRC4 %V([14]) filesrc4
.model filesrc4 filesource (file="dat/y2_profile_bunched.txt" amploffset=[0 0] amplscale=[1 1]
+ timeoffset=0 timescale=1
+ timerelative=false amplstep=false) )

.CONTROL

TRAN 20ns 4ms
*AC DEC 5 10 1000MEG 
plot v(1) v(2)
plot v(11) v(22)
plot v(13) v(23)
plot v(14) v(24)
wrdata x1_bunched_100k_20ns (V(2))
wrdata x2_bunched_100k_20ns (V(22)) 
wrdata y1_bunched_100k_20ns (V(23)) 
wrdata y2_bunched_100k_20ns (V(24)) 

*wrdata mag50 (v(22)) 
*wrdata magnitude1 (V(2)) 
*wrdata phase1 phase(v(2)) 
*wrdata magnitude2 (V(23)) 
*wrdata phase2 phase(v(23))
*wrdata magnitude3 (V(22)) 
*wrdata phase3 phase(v(22))  
*.include freq_analysis.txt
*.include plotng.txt

.endc
.END

  
