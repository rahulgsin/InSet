* Version 2.0 Copyright © Linear Technology Corp. 10/19/05. All rights reserved.
*
.SUBCKT LT1363 3 2 7 4 6 ;(+IN -IN V+ V- OUT)
* INPUT
RC1 7 80 568.41
RC2 7 90 568.41
Q1 80 2 10 QM1
Q2 90 3 11 QM2
CIN 2 3 2e-12
*INPUT POLE AT 300MHZ
C1 80 90 4.67e-13
RE1 10 12 555.32
RE2 11 12 555.32
IEE 12 4 0.0040012
RE 12 0 49985
* INTERMEDIATE
GCM 8 0 12 0 5.5634e-8
GA 8 0 78 0 0.0017593
R2 8 0 3690000
C2 8 0 3.85E-12
DC1 8 7 DM3
DC2 4 8 DM3
*
*POLE AT 300MHZ
GX1 0 28 90 80 1E-06
RX1 28 0 1E+06
CX1 28 0 5.3e-16
*POLE AT 300MHZ
GX2 0 38 28 0 1E-06
RX2 38 0 1E+06
CX2 38 0 5.3e-16
*POLE AT 300MHZ
GX3 0 48 38 0 1E-06
RX3 48 0 1E+06
CX3 48 0 5.3e-16
*ZERO AT 85MHZ
GX4 0 58 48 0 1E-06
RX4 58 59 1E+06
LX4 59 0 0.00187
*POLE AT 170MHZ
GX5 0 68 58 0 1E-06
RX5 68 0 1E+06
CX5 68 0 9.37e-16
*POLE AT 500MHZ
GX6 0 78 68 0 1E-06
RX6 78 0 1E+06
CX6 78 0 3.18e-16
*
EB 1 0 8 0 1
RO2 1 6 20
RF 8 99 800
CF 99 6 6E-12
* OUTPUT
ECL 18 1 6 1 0.36
Q3 7 18 8 QM3
Q4 4 18 8 QM4
*
D3A 131 70 DM3
D3B 13 131 DM3
GPL 8 0 70 7 1
VC 13 6 2.9317
RPLA 7 70 10
RPLB 7 131 1000
D4A 60 141 DM3
D4B 141 14 DM3
GNL 8 0 60 4 1
VE 6 14 2.9317
RNLA 60 4 10
RNLB 141 4 1000
*
IP 7 4 0.0019988
DSUB 4 7 DM2
* MODELS
.MODEL QM1 NPN(IS=8e-16 BF=3030.3)
.MODEL QM2 NPN(IS=8.1562E-16 BF=3703.7)
.MODEL QM3 NPN(IS=8e-16 BF=100)
.MODEL QM4 PNP(IS=8e-16 BF=100)
.MODEL DM1 D(IS=1e-20)
.MODEL DM2 D(IS=8e-16 BV=43.2)
.MODEL DM3 D(IS=1e-16)
.ENDS LT1363
*

